library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity program_counter is

end entity program_counter;

architecture Behavior of program_counter is

end architecture Behavior;

